XlxV38EB    1173     5df�%<��z�N�Eh��%b��!I;YcB=p������$AH[v���"E{8$�\$2d���5����53/%!�4��3�6zo-��Bfa��G^�^�JL����x�:�����O��&�-*�/���f'��z	����J���Z4@a&FN'h���k��)��r�$O) �#�Z>:H�.+�*�*�Z!���̊��I�UxI�A�϶$T���������a����g���C BwN�����e"�����������n�<E�$S�v�!�W�%�D�)͂�J ��cl��dW���)5Z�	�cS'+6�0�TY� �@˘}�a�Z
}]S�m���4��xn�5��$����G���<c�Ŕ��|�+{f��\N*J�rb���-`
P2z���aN�0a�}��y�4��P=d�B3���+RK��U�a����&��~Y�g��:t��#�	�v���^a 〘� a� �r�2�s}_�E�1�h�� �Y��&V�O�x��<��f��� �Q�ߧ��YƸK����>����l>�,�ܫ�~:r^��	�s!��R��c3�B�%z��R'�nHt�vZ��U�N��U4�PD��h�K��,=��-0�fp$h�����XH�[�ZuW8��NͿ@� dD�1�W�`f'y��ҟ��@��4�]�(�M/ b����К��V�_G�CsGF6�{�5C+/�aFR�9%��vD��!s���5^�	0��Vԭ�tn����@ۉ(d���"R�,:gt��!��s#Q�����<��"�_S/�@��|߹D�as���6L(~n-��e )}aWh401������|��7���y{��n�� m�r�B�:�f_$\���p��ڲ|ԉP��EXgQ�>ᶡ�8;^� ���Q��'I�Q��ˈXR��#�>�"H��P-�ݼ�*�7b����ƾb�N������|R��'��J:<@`��ܮzޅA�O���OGD@p�7š5�/�=P���B�h��T��Z�B�ˇ�d$�8\�魡�W�V��/�:�*��9^�nI�� ��DA<uN9�fl���%L�fm_�Zn�Ƙa�m'K���rC�ǌ��u�O��u�܁�-�t��#�9�_�����oe�;N����4^%�	C���9�* � O厫┡�o�@e�6wj_C>s!&:�g{��݅
��N���+�95�x0Ȯ`�g��|���n� Y��z������V+�t�y_��#}�A�ⴷ�u�9����#R��z� >1G�sMP	�}s�a�i���r�_��N�*��=?L2��	�,���p�%ưSf�����E���B�g��}I������k�چ��������jo�(�~�K�ș�g�|�ǚ�� k$9���d��V�[O�l~4��¿5h����5 �������Y��'��K9�����J~`����<�Z9?:<�aZBbS� C��