XlxV38EB    109c     5d6�uW
��*v�Ifɽ�^Ƅ�����L�[��sp�NvdB��@�y?IG��b\���ӱ����ۡ�q��$^h�Cb�a�?Z뇮�q9���s�,�ŀ|�613�C�PQ������K�U����c��ޯ��v�]�Hnh��;}��W��j�.�-��UHx**{�씀�ׯG��uqe���D�i�ː�����E�#�Ri/�è
�Mo�o�r�� &�{�>�O{9��Gf�݌[�Jf�Nn�.���&��žk��>d�(����n=\i�Lm��C�N;Q�S�}y��un���Q����OYLx�[��{k춳׶��ҮHS5D�_�y�����g-�""��R5o]�x�iS�M����%!��iܭ�TĢ�ɶ;j��!x���N���>������� ��y1�]�)wt���|���sX�}ƹ$� �ɧ@�2}�@�-���k�n�?c�V�0��A[��� ���z��>K�n��Dn�E�L%�����ǉ�P��u������X��
��E5='��Pa��'��+�L���/�U�KfF �xo[�~�қ�M3�r�$w�n1���v�Wƚ�1�ݒ@��u>�=��;�o��O�Ku(��?���Q"�,���,�Ǣ��t��T�h̋��p{����,'�	V�d��%����:?����Չ�h���acj� �̚�@7��\�|5�wR�M�2!�x�;8��/g����U��)��g��t?T�����{5ߵj;o��A��[A��t�J���6�v�B�m?��H��pԲ1�{�;r�sD���M7�ߋm��b����'�O���+#SlS�f#ZVa���mf�T�(6�ow��E��|R�_��}�����'���Tꗗ]�ܩ�_�ڻ��a���]�~�q��M(<ߘ� _`���7Vǡ��ؾ�3��	F`�'V��]7O$�8_GZ���([ާ�9��'�h�����p����&��r�H���Z?��U�����Uv�#�k�ɘ#$Gm�!�c����P���	�k�K�:����D���|f!���׿�P֍"Y�<q1a��|��맲�'��J\�K��;t-<¡�6^>��[���W���$|{w|'�R�������Y8�Ȁ�����x��Ek����e�Q�$O���=.������i0��_�d}]:nW̤e���X���U�����޴�h��K�}v)
��c�I�d���{���Z��j�A�6��l��)� 1tﯠ�O�(U�TQ�3����8�X����>)'1�IKM�*xٺ�R_I��w�7�r�*�r��N���U�>�;�W��HIA�s9]����2!T��t�N�R%�/�~��oJ4t����l}�5�E�8;�\�D6��O��������M�jY��s�$Iu�V���ט�I8`?��?���=��h�^}wu�n:H9�e����H)N ��}